magic
tech scmos
magscale 1 2
timestamp 1600036315
<< metal1 >>
rect 474 814 486 816
rect 459 806 461 814
rect 469 806 471 814
rect 479 806 481 814
rect 489 806 491 814
rect 499 806 501 814
rect 474 804 486 806
rect 100 697 131 703
rect 540 697 563 703
rect 540 692 548 697
rect 970 614 982 616
rect 955 606 957 614
rect 965 606 967 614
rect 975 606 977 614
rect 985 606 987 614
rect 995 606 997 614
rect 970 604 982 606
rect 728 537 748 543
rect 957 537 1020 543
rect 173 517 211 523
rect 221 517 259 523
rect 301 503 307 528
rect 541 517 572 523
rect 900 517 915 523
rect 316 512 324 516
rect 301 497 323 503
rect 340 497 356 503
rect 348 492 356 497
rect 669 497 684 503
rect 474 414 486 416
rect 459 406 461 414
rect 469 406 471 414
rect 479 406 481 414
rect 489 406 491 414
rect 499 406 501 414
rect 474 404 486 406
rect 93 317 108 323
rect 877 317 892 323
rect 125 297 140 303
rect 157 297 195 303
rect 317 297 332 303
rect 516 277 547 283
rect 573 283 579 303
rect 573 277 652 283
rect 941 277 956 283
rect 84 256 92 264
rect 420 257 435 263
rect 628 257 659 263
rect 970 214 982 216
rect 955 206 957 214
rect 965 206 967 214
rect 975 206 977 214
rect 985 206 987 214
rect 995 206 997 214
rect 970 204 982 206
rect 522 176 524 184
rect 188 137 212 143
rect 589 117 612 123
rect 604 114 612 117
rect 474 14 486 16
rect 459 6 461 14
rect 469 6 471 14
rect 479 6 481 14
rect 489 6 491 14
rect 499 6 501 14
rect 474 4 486 6
<< m2contact >>
rect 451 806 459 814
rect 461 806 469 814
rect 471 806 479 814
rect 481 806 489 814
rect 491 806 499 814
rect 501 806 509 814
rect 236 776 244 784
rect 444 776 452 784
rect 588 776 596 784
rect 92 696 100 704
rect 204 696 212 704
rect 300 694 308 702
rect 476 696 484 704
rect 524 696 532 704
rect 716 696 724 704
rect 908 696 916 704
rect 172 676 180 684
rect 332 676 340 684
rect 540 676 548 684
rect 716 676 724 684
rect 764 676 772 684
rect 892 676 900 684
rect 12 636 20 644
rect 428 636 436 644
rect 492 636 500 644
rect 604 636 612 644
rect 796 636 804 644
rect 947 606 955 614
rect 957 606 965 614
rect 967 606 975 614
rect 977 606 985 614
rect 987 606 995 614
rect 997 606 1005 614
rect 44 576 52 584
rect 156 576 164 584
rect 252 576 260 584
rect 588 576 596 584
rect 812 576 820 584
rect 844 576 852 584
rect 60 556 68 564
rect 140 556 148 564
rect 572 556 580 564
rect 684 556 692 564
rect 828 556 836 564
rect 28 536 36 544
rect 76 536 84 544
rect 108 536 116 544
rect 236 536 244 544
rect 380 536 388 544
rect 460 536 468 544
rect 508 536 516 544
rect 620 536 628 544
rect 668 536 676 544
rect 748 536 756 544
rect 796 536 804 544
rect 892 536 900 544
rect 1020 536 1028 544
rect 12 516 20 524
rect 92 516 100 524
rect 284 516 292 524
rect 124 496 132 504
rect 188 496 196 504
rect 316 516 324 524
rect 332 516 340 524
rect 396 516 404 524
rect 476 516 484 524
rect 524 516 532 524
rect 572 516 580 524
rect 604 516 612 524
rect 636 516 644 524
rect 748 516 756 524
rect 780 516 788 524
rect 876 516 884 524
rect 892 516 900 524
rect 924 516 932 524
rect 332 496 340 504
rect 428 496 436 504
rect 492 496 500 504
rect 556 496 564 504
rect 684 496 692 504
rect 700 496 708 504
rect 764 496 772 504
rect 460 476 468 484
rect 732 476 740 484
rect 332 436 340 444
rect 451 406 459 414
rect 461 406 469 414
rect 471 406 479 414
rect 481 406 489 414
rect 491 406 499 414
rect 501 406 509 414
rect 732 376 740 384
rect 108 316 116 324
rect 172 316 180 324
rect 252 316 260 324
rect 284 316 292 324
rect 348 316 356 324
rect 460 316 468 324
rect 892 316 900 324
rect 44 296 52 304
rect 140 296 148 304
rect 332 296 340 304
rect 380 296 388 304
rect 412 296 420 304
rect 12 276 20 284
rect 60 276 68 284
rect 140 276 148 284
rect 204 276 212 284
rect 268 276 276 284
rect 284 276 292 284
rect 332 276 340 284
rect 364 276 372 284
rect 396 276 404 284
rect 492 276 500 284
rect 508 276 516 284
rect 556 276 564 284
rect 588 296 596 304
rect 684 296 692 304
rect 764 296 772 304
rect 844 296 852 304
rect 924 296 932 304
rect 1004 296 1012 304
rect 652 276 660 284
rect 668 276 676 284
rect 780 276 788 284
rect 828 276 836 284
rect 860 276 868 284
rect 908 276 916 284
rect 956 276 964 284
rect 988 276 996 284
rect 92 256 100 264
rect 108 256 116 264
rect 236 256 244 264
rect 412 256 420 264
rect 444 256 452 264
rect 508 256 516 264
rect 524 256 532 264
rect 620 256 628 264
rect 812 256 820 264
rect 956 256 964 264
rect 220 236 228 244
rect 796 236 804 244
rect 972 236 980 244
rect 947 206 955 214
rect 957 206 965 214
rect 967 206 975 214
rect 977 206 985 214
rect 987 206 995 214
rect 997 206 1005 214
rect 12 176 20 184
rect 444 176 452 184
rect 524 176 532 184
rect 604 176 612 184
rect 796 176 804 184
rect 492 136 500 144
rect 540 136 548 144
rect 716 136 724 144
rect 140 118 148 126
rect 268 116 276 124
rect 316 116 324 124
rect 428 116 436 124
rect 476 116 484 124
rect 732 118 740 126
rect 860 116 868 124
rect 924 118 932 126
rect 508 96 516 104
rect 380 76 388 84
rect 396 36 404 44
rect 556 36 564 44
rect 451 6 459 14
rect 461 6 469 14
rect 471 6 479 14
rect 481 6 489 14
rect 491 6 499 14
rect 501 6 509 14
<< metal2 >>
rect 221 857 243 863
rect 237 784 243 857
rect 474 814 486 816
rect 459 806 461 814
rect 469 806 471 814
rect 479 806 481 814
rect 489 806 491 814
rect 499 806 501 814
rect 474 804 486 806
rect 541 784 547 863
rect 13 644 19 696
rect 93 684 99 696
rect 13 524 19 636
rect 45 584 51 676
rect 301 624 307 694
rect 429 644 435 696
rect 157 584 163 616
rect 429 603 435 636
rect 413 597 435 603
rect 253 564 259 576
rect 61 544 67 556
rect 29 504 35 536
rect 77 524 83 536
rect 141 524 147 556
rect 13 284 19 296
rect 45 184 51 296
rect 61 284 67 516
rect 125 444 131 496
rect 141 324 147 516
rect 237 504 243 536
rect 317 524 323 536
rect 333 524 339 576
rect 189 444 195 496
rect 397 464 403 516
rect 413 504 419 597
rect 461 524 467 536
rect 461 484 467 496
rect 477 484 483 516
rect 493 504 499 636
rect 509 544 515 616
rect 541 583 547 676
rect 573 624 579 863
rect 589 857 611 863
rect 589 784 595 857
rect 589 584 595 696
rect 605 584 611 636
rect 532 577 547 583
rect 525 524 531 576
rect 685 564 691 636
rect 557 484 563 496
rect 109 304 115 316
rect 333 304 339 436
rect 349 324 355 436
rect 381 304 387 316
rect 109 264 115 296
rect 205 284 211 296
rect 269 284 275 296
rect 397 284 403 296
rect 413 284 419 296
rect 237 264 243 276
rect 333 264 339 276
rect 221 124 227 236
rect 413 164 419 256
rect 429 243 435 476
rect 557 444 563 476
rect 474 414 486 416
rect 459 406 461 414
rect 469 406 471 414
rect 479 406 481 414
rect 489 406 491 414
rect 499 406 501 414
rect 474 404 486 406
rect 445 264 451 276
rect 493 244 499 276
rect 429 237 451 243
rect 445 184 451 237
rect 493 184 499 236
rect 525 203 531 256
rect 509 197 531 203
rect 269 124 275 156
rect 493 144 499 156
rect 317 124 323 136
rect 509 124 515 197
rect 557 184 563 276
rect 621 264 627 536
rect 637 524 643 536
rect 669 524 675 536
rect 685 504 691 556
rect 669 244 675 276
rect 541 164 547 176
rect 541 144 547 156
rect 717 144 723 676
rect 813 584 819 696
rect 861 623 867 863
rect 845 617 867 623
rect 845 584 851 617
rect 877 524 883 636
rect 970 614 982 616
rect 955 606 957 614
rect 965 606 967 614
rect 975 606 977 614
rect 985 606 987 614
rect 995 606 997 614
rect 970 604 982 606
rect 893 544 899 556
rect 1021 524 1027 536
rect 749 504 755 516
rect 733 384 739 476
rect 765 464 771 496
rect 893 484 899 516
rect 765 404 771 456
rect 733 304 739 376
rect 893 324 899 476
rect 925 404 931 516
rect 765 244 771 296
rect 845 284 851 296
rect 957 284 963 396
rect 989 284 995 296
rect 1005 284 1011 296
rect 829 244 835 276
rect 861 264 867 276
rect 909 264 915 276
rect 765 184 771 236
rect 797 203 803 236
rect 797 197 819 203
rect 813 124 819 197
rect 861 124 867 136
rect 925 126 931 236
rect 970 214 982 216
rect 955 206 957 214
rect 965 206 967 214
rect 975 206 977 214
rect 985 206 987 214
rect 995 206 997 214
rect 970 204 982 206
rect 381 84 387 116
rect 509 104 515 116
rect 397 -17 403 36
rect 474 14 486 16
rect 459 6 461 14
rect 469 6 471 14
rect 479 6 481 14
rect 489 6 491 14
rect 499 6 501 14
rect 474 4 486 6
rect 557 -17 563 36
rect 397 -23 419 -17
rect 557 -23 579 -17
<< m3contact >>
rect 451 806 459 814
rect 461 806 469 814
rect 471 806 479 814
rect 481 806 489 814
rect 491 806 499 814
rect 501 806 509 814
rect 444 776 452 784
rect 540 776 548 784
rect 12 696 20 704
rect 204 696 212 704
rect 428 696 436 704
rect 476 696 484 704
rect 524 696 532 704
rect 44 676 52 684
rect 92 676 100 684
rect 172 676 180 684
rect 332 676 340 684
rect 156 616 164 624
rect 300 616 308 624
rect 332 576 340 584
rect 252 556 260 564
rect 60 536 68 544
rect 108 536 116 544
rect 12 516 20 524
rect 316 536 324 544
rect 60 516 68 524
rect 76 516 84 524
rect 92 516 100 524
rect 140 516 148 524
rect 28 496 36 504
rect 12 296 20 304
rect 44 296 52 304
rect 124 436 132 444
rect 380 536 388 544
rect 284 516 292 524
rect 332 516 340 524
rect 236 496 244 504
rect 332 496 340 504
rect 460 516 468 524
rect 412 496 420 504
rect 428 496 436 504
rect 460 496 468 504
rect 508 616 516 624
rect 524 576 532 584
rect 588 696 596 704
rect 716 696 724 704
rect 812 696 820 704
rect 572 616 580 624
rect 764 676 772 684
rect 684 636 692 644
rect 604 576 612 584
rect 508 536 516 544
rect 572 556 580 564
rect 636 536 644 544
rect 572 516 580 524
rect 604 516 612 524
rect 428 476 436 484
rect 476 476 484 484
rect 556 476 564 484
rect 396 456 404 464
rect 188 436 196 444
rect 348 436 356 444
rect 140 316 148 324
rect 172 316 180 324
rect 252 316 260 324
rect 284 316 292 324
rect 348 316 356 324
rect 380 316 388 324
rect 108 296 116 304
rect 140 296 148 304
rect 204 296 212 304
rect 268 296 276 304
rect 332 296 340 304
rect 396 296 404 304
rect 60 276 68 284
rect 140 276 148 284
rect 236 276 244 284
rect 284 276 292 284
rect 364 276 372 284
rect 412 276 420 284
rect 92 256 100 264
rect 332 256 340 264
rect 12 176 20 184
rect 44 176 52 184
rect 556 436 564 444
rect 451 406 459 414
rect 461 406 469 414
rect 471 406 479 414
rect 481 406 489 414
rect 491 406 499 414
rect 501 406 509 414
rect 460 316 468 324
rect 588 296 596 304
rect 444 276 452 284
rect 508 276 516 284
rect 508 256 516 264
rect 492 236 500 244
rect 492 176 500 184
rect 268 156 276 164
rect 412 156 420 164
rect 492 156 500 164
rect 316 136 324 144
rect 668 516 676 524
rect 700 496 708 504
rect 684 296 692 304
rect 652 276 660 284
rect 620 256 628 264
rect 668 236 676 244
rect 524 176 532 184
rect 540 176 548 184
rect 556 176 564 184
rect 604 176 612 184
rect 540 156 548 164
rect 796 636 804 644
rect 908 696 916 704
rect 892 676 900 684
rect 876 636 884 644
rect 828 556 836 564
rect 748 536 756 544
rect 796 536 804 544
rect 947 606 955 614
rect 957 606 965 614
rect 967 606 975 614
rect 977 606 985 614
rect 987 606 995 614
rect 997 606 1005 614
rect 892 556 900 564
rect 780 516 788 524
rect 1020 516 1028 524
rect 748 496 756 504
rect 892 476 900 484
rect 764 456 772 464
rect 764 396 772 404
rect 924 396 932 404
rect 956 396 964 404
rect 732 296 740 304
rect 924 296 932 304
rect 988 296 996 304
rect 780 276 788 284
rect 844 276 852 284
rect 956 276 964 284
rect 1004 276 1012 284
rect 812 256 820 264
rect 860 256 868 264
rect 908 256 916 264
rect 956 256 964 264
rect 764 236 772 244
rect 828 236 836 244
rect 924 236 932 244
rect 972 236 980 244
rect 764 176 772 184
rect 796 176 804 184
rect 716 136 724 144
rect 860 136 868 144
rect 947 206 955 214
rect 957 206 965 214
rect 967 206 975 214
rect 977 206 985 214
rect 987 206 995 214
rect 997 206 1005 214
rect 140 118 148 124
rect 140 116 148 118
rect 220 116 228 124
rect 380 116 388 124
rect 428 116 436 124
rect 476 116 484 124
rect 508 116 516 124
rect 732 118 740 124
rect 732 116 740 118
rect 812 116 820 124
rect 451 6 459 14
rect 461 6 469 14
rect 471 6 479 14
rect 481 6 489 14
rect 491 6 499 14
rect 501 6 509 14
<< metal3 >>
rect 450 814 510 816
rect 450 806 451 814
rect 460 806 461 814
rect 499 806 500 814
rect 509 806 510 814
rect 450 804 510 806
rect 452 777 540 783
rect 20 697 204 703
rect 436 697 476 703
rect 484 697 524 703
rect 596 697 716 703
rect 820 697 908 703
rect 52 677 92 683
rect 180 677 332 683
rect 340 677 764 683
rect 772 677 892 683
rect 900 677 1059 683
rect 692 637 796 643
rect 804 637 876 643
rect 164 617 300 623
rect 516 617 572 623
rect 946 614 1006 616
rect 946 606 947 614
rect 956 606 957 614
rect 995 606 996 614
rect 1005 606 1006 614
rect 946 604 1006 606
rect 340 577 524 583
rect 532 577 604 583
rect 260 557 572 563
rect 836 557 892 563
rect 900 557 1059 563
rect 68 537 108 543
rect 324 537 380 543
rect 388 537 508 543
rect 557 537 636 543
rect 20 517 60 523
rect 68 517 76 523
rect 100 517 140 523
rect 292 517 332 523
rect 557 523 563 537
rect 756 537 796 543
rect 468 517 563 523
rect 580 517 604 523
rect 676 517 780 523
rect 1028 517 1059 523
rect 93 503 99 516
rect 36 497 99 503
rect 244 497 332 503
rect 340 497 412 503
rect 436 497 460 503
rect 708 497 748 503
rect 436 477 476 483
rect 564 477 892 483
rect 404 457 764 463
rect 132 437 188 443
rect 196 437 348 443
rect 356 437 556 443
rect 450 414 510 416
rect 450 406 451 414
rect 460 406 461 414
rect 499 406 500 414
rect 509 406 510 414
rect 450 404 510 406
rect 772 397 780 403
rect 788 397 924 403
rect 932 397 956 403
rect 148 317 172 323
rect 180 317 252 323
rect 292 317 348 323
rect 388 317 460 323
rect -35 297 12 303
rect 52 297 108 303
rect 148 297 204 303
rect 276 297 332 303
rect 340 297 396 303
rect 404 297 588 303
rect 596 297 684 303
rect 740 297 924 303
rect 932 297 988 303
rect 68 277 140 283
rect 244 277 284 283
rect 372 277 412 283
rect 452 277 508 283
rect 660 277 780 283
rect 788 277 844 283
rect 964 277 1004 283
rect 100 257 332 263
rect 340 257 508 263
rect 516 257 620 263
rect 820 257 860 263
rect 916 257 956 263
rect 500 237 668 243
rect 772 237 828 243
rect 932 237 972 243
rect 946 214 1006 216
rect 946 206 947 214
rect 956 206 957 214
rect 995 206 996 214
rect 1005 206 1006 214
rect 946 204 1006 206
rect 20 177 44 183
rect 500 177 524 183
rect 548 177 556 183
rect 564 177 604 183
rect 612 177 764 183
rect 788 177 796 183
rect 276 157 412 163
rect 500 157 540 163
rect 324 137 716 143
rect 724 137 860 143
rect 148 117 220 123
rect 388 117 428 123
rect 436 117 476 123
rect 484 117 508 123
rect 740 117 812 123
rect 450 14 510 16
rect 450 6 451 14
rect 460 6 461 14
rect 499 6 500 14
rect 509 6 510 14
rect 450 4 510 6
<< m4contact >>
rect 452 806 459 814
rect 459 806 460 814
rect 464 806 469 814
rect 469 806 471 814
rect 471 806 472 814
rect 476 806 479 814
rect 479 806 481 814
rect 481 806 484 814
rect 488 806 489 814
rect 489 806 491 814
rect 491 806 496 814
rect 500 806 501 814
rect 501 806 508 814
rect 948 606 955 614
rect 955 606 956 614
rect 960 606 965 614
rect 965 606 967 614
rect 967 606 968 614
rect 972 606 975 614
rect 975 606 977 614
rect 977 606 980 614
rect 984 606 985 614
rect 985 606 987 614
rect 987 606 992 614
rect 996 606 997 614
rect 997 606 1004 614
rect 452 406 459 414
rect 459 406 460 414
rect 464 406 469 414
rect 469 406 471 414
rect 471 406 472 414
rect 476 406 479 414
rect 479 406 481 414
rect 481 406 484 414
rect 488 406 489 414
rect 489 406 491 414
rect 491 406 496 414
rect 500 406 501 414
rect 501 406 508 414
rect 780 396 788 404
rect 948 206 955 214
rect 955 206 956 214
rect 960 206 965 214
rect 965 206 967 214
rect 967 206 968 214
rect 972 206 975 214
rect 975 206 977 214
rect 977 206 980 214
rect 984 206 985 214
rect 985 206 987 214
rect 987 206 992 214
rect 996 206 997 214
rect 997 206 1004 214
rect 780 176 788 184
rect 452 6 459 14
rect 459 6 460 14
rect 464 6 469 14
rect 469 6 471 14
rect 471 6 472 14
rect 476 6 479 14
rect 479 6 481 14
rect 481 6 484 14
rect 488 6 489 14
rect 489 6 491 14
rect 491 6 496 14
rect 500 6 501 14
rect 501 6 508 14
<< metal4 >>
rect 448 814 512 816
rect 448 806 452 814
rect 460 806 464 814
rect 472 806 476 814
rect 484 806 488 814
rect 496 806 500 814
rect 508 806 512 814
rect 448 414 512 806
rect 448 406 452 414
rect 460 406 464 414
rect 472 406 476 414
rect 484 406 488 414
rect 496 406 500 414
rect 508 406 512 414
rect 944 614 1008 816
rect 944 606 948 614
rect 956 606 960 614
rect 968 606 972 614
rect 980 606 984 614
rect 992 606 996 614
rect 1004 606 1008 614
rect 448 14 512 406
rect 778 404 790 406
rect 778 396 780 404
rect 788 396 790 404
rect 778 184 790 396
rect 778 176 780 184
rect 788 176 790 184
rect 778 174 790 176
rect 944 214 1008 606
rect 944 206 948 214
rect 956 206 960 214
rect 968 206 972 214
rect 980 206 984 214
rect 992 206 996 214
rect 1004 206 1008 214
rect 448 6 452 14
rect 460 6 464 14
rect 472 6 476 14
rect 484 6 488 14
rect 496 6 500 14
rect 508 6 512 14
rect 448 -10 512 6
rect 944 -10 1008 206
use DFFPOSX1  _73_
timestamp 1600036315
transform -1 0 200 0 -1 210
box -4 -6 196 206
use DFFPOSX1  _75_
timestamp 1600036315
transform 1 0 200 0 -1 210
box -4 -6 196 206
use BUFX2  _65_
timestamp 1600036315
transform -1 0 56 0 1 210
box -4 -6 52 206
use NAND2X1  _40_
timestamp 1600036315
transform 1 0 56 0 1 210
box -4 -6 52 206
use INVX1  _38_
timestamp 1600036315
transform 1 0 104 0 1 210
box -4 -6 36 206
use NAND2X1  _39_
timestamp 1600036315
transform 1 0 136 0 1 210
box -4 -6 52 206
use AOI21X1  _42_
timestamp 1600036315
transform 1 0 184 0 1 210
box -4 -6 68 206
use BUFX2  _67_
timestamp 1600036315
transform -1 0 440 0 -1 210
box -4 -6 52 206
use INVX2  _33_
timestamp 1600036315
transform -1 0 280 0 1 210
box -4 -6 36 206
use OAI21X1  _41_
timestamp 1600036315
transform -1 0 344 0 1 210
box -4 -6 68 206
use OAI21X1  _49_
timestamp 1600036315
transform -1 0 408 0 1 210
box -4 -6 68 206
use NOR2X1  _50_
timestamp 1600036315
transform -1 0 456 0 1 210
box -4 -6 52 206
use AND2X2  _55_
timestamp 1600036315
transform -1 0 504 0 -1 210
box -4 -6 68 206
use NAND2X1  _47_
timestamp 1600036315
transform -1 0 552 0 -1 210
box -4 -6 52 206
use BUFX2  _66_
timestamp 1600036315
transform -1 0 600 0 -1 210
box -4 -6 52 206
use DFFPOSX1  _74_
timestamp 1600036315
transform -1 0 792 0 -1 210
box -4 -6 196 206
use OR2X2  _48_
timestamp 1600036315
transform -1 0 520 0 1 210
box -4 -6 68 206
use AOI21X1  _46_
timestamp 1600036315
transform -1 0 584 0 1 210
box -4 -6 68 206
use NOR2X1  _43_
timestamp 1600036315
transform -1 0 632 0 1 210
box -4 -6 52 206
use DFFPOSX1  _76_
timestamp 1600036315
transform -1 0 984 0 -1 210
box -4 -6 196 206
use NOR3X1  _51_
timestamp 1600036315
transform 1 0 632 0 1 210
box -4 -6 132 206
use AOI21X1  _45_
timestamp 1600036315
transform 1 0 760 0 1 210
box -4 -6 68 206
use OAI21X1  _44_
timestamp 1600036315
transform 1 0 824 0 1 210
box -4 -6 68 206
use OAI21X1  _52_
timestamp 1600036315
transform -1 0 952 0 1 210
box -4 -6 68 206
use AOI21X1  _53_
timestamp 1600036315
transform -1 0 1016 0 1 210
box -4 -6 68 206
use FILL  FILL9840x100
timestamp 1600036315
transform -1 0 1000 0 -1 210
box -4 -6 20 206
use FILL  FILL10000x100
timestamp 1600036315
transform -1 0 1016 0 -1 210
box -4 -6 20 206
use AOI21X1  _37_
timestamp 1600036315
transform 1 0 8 0 -1 610
box -4 -6 68 206
use OAI21X1  _36_
timestamp 1600036315
transform 1 0 72 0 -1 610
box -4 -6 68 206
use NOR2X1  _35_
timestamp 1600036315
transform 1 0 136 0 -1 610
box -4 -6 52 206
use OAI21X1  _34_
timestamp 1600036315
transform -1 0 248 0 -1 610
box -4 -6 68 206
use AND2X2  _28_
timestamp 1600036315
transform -1 0 312 0 -1 610
box -4 -6 68 206
use NAND3X1  _32_
timestamp 1600036315
transform 1 0 312 0 -1 610
box -4 -6 68 206
use AND2X2  _56_
timestamp 1600036315
transform 1 0 376 0 -1 610
box -4 -6 68 206
use NAND3X1  _57_
timestamp 1600036315
transform -1 0 504 0 -1 610
box -4 -6 68 206
use OAI21X1  _30_
timestamp 1600036315
transform 1 0 504 0 -1 610
box -4 -6 68 206
use NOR2X1  _31_
timestamp 1600036315
transform 1 0 568 0 -1 610
box -4 -6 52 206
use OAI21X1  _58_
timestamp 1600036315
transform 1 0 616 0 -1 610
box -4 -6 68 206
use INVX1  _59_
timestamp 1600036315
transform 1 0 680 0 -1 610
box -4 -6 36 206
use NAND3X1  _60_
timestamp 1600036315
transform -1 0 776 0 -1 610
box -4 -6 68 206
use AOI21X1  _61_
timestamp 1600036315
transform 1 0 776 0 -1 610
box -4 -6 68 206
use BUFX2  _69_
timestamp 1600036315
transform -1 0 888 0 -1 610
box -4 -6 52 206
use INVX2  _29_
timestamp 1600036315
transform 1 0 888 0 -1 610
box -4 -6 36 206
use BUFX2  _68_
timestamp 1600036315
transform 1 0 920 0 -1 610
box -4 -6 52 206
use FILL  FILL9680x4100
timestamp 1600036315
transform -1 0 984 0 -1 610
box -4 -6 20 206
use FILL  FILL9840x4100
timestamp 1600036315
transform -1 0 1000 0 -1 610
box -4 -6 20 206
use FILL  FILL10000x4100
timestamp 1600036315
transform -1 0 1016 0 -1 610
box -4 -6 20 206
use DFFPOSX1  _72_
timestamp 1600036315
transform -1 0 200 0 1 610
box -4 -6 196 206
use BUFX2  _64_
timestamp 1600036315
transform 1 0 200 0 1 610
box -4 -6 52 206
use DFFPOSX1  _71_
timestamp 1600036315
transform 1 0 248 0 1 610
box -4 -6 196 206
use BUFX2  _63_
timestamp 1600036315
transform -1 0 488 0 1 610
box -4 -6 52 206
use AND2X2  _54_
timestamp 1600036315
transform -1 0 552 0 1 610
box -4 -6 68 206
use BUFX2  _62_
timestamp 1600036315
transform 1 0 552 0 1 610
box -4 -6 52 206
use DFFPOSX1  _70_
timestamp 1600036315
transform -1 0 792 0 1 610
box -4 -6 196 206
use DFFPOSX1  _77_
timestamp 1600036315
transform -1 0 984 0 1 610
box -4 -6 196 206
use FILL  FILL9840x6100
timestamp 1600036315
transform 1 0 984 0 1 610
box -4 -6 20 206
use FILL  FILL10000x6100
timestamp 1600036315
transform 1 0 1000 0 1 610
box -4 -6 20 206
<< labels >>
rlabel metal4 s 944 -10 1008 0 8 gnd
port 0 nsew
rlabel metal4 s 448 -10 512 0 8 vdd
port 1 nsew
rlabel metal3 s 1053 677 1059 683 6 clk
port 2 nsew
rlabel metal2 s 861 857 867 863 6 count[7]
port 3 nsew
rlabel metal3 s 1053 517 1059 523 6 count[6]
port 4 nsew
rlabel metal2 s 413 -23 419 -17 8 count[5]
port 5 nsew
rlabel metal2 s 573 -23 579 -17 8 count[4]
port 6 nsew
rlabel metal3 s -35 297 -29 303 4 count[3]
port 7 nsew
rlabel metal2 s 221 857 227 863 6 count[2]
port 8 nsew
rlabel metal2 s 541 857 547 863 6 count[1]
port 9 nsew
rlabel metal2 s 605 857 611 863 6 count[0]
port 10 nsew
rlabel metal2 s 573 857 579 863 6 en
port 11 nsew
rlabel metal3 s 1053 557 1059 563 6 rst
port 12 nsew
<< end >>
