magic
tech scmos
magscale 1 2
timestamp 1600036665
<< checkpaint >>
rect -76 -66 140 270
<< nwell >>
rect -16 96 80 210
<< ntransistor >>
rect 14 12 18 52
rect 24 12 28 52
rect 40 12 44 52
<< ptransistor >>
rect 14 148 18 188
rect 30 148 34 188
rect 46 108 50 188
<< ndiffusion >>
rect 4 51 14 52
rect 12 13 14 51
rect 4 12 14 13
rect 18 12 24 52
rect 28 50 40 52
rect 28 12 30 50
rect 38 12 40 50
rect 44 51 54 52
rect 44 13 46 51
rect 44 12 54 13
<< pdiffusion >>
rect 4 187 14 188
rect 12 149 14 187
rect 4 148 14 149
rect 18 187 30 188
rect 18 149 20 187
rect 28 149 30 187
rect 18 148 30 149
rect 34 184 46 188
rect 34 148 36 184
rect 44 116 46 184
rect 36 112 46 116
rect 40 108 46 112
rect 50 187 60 188
rect 50 109 52 187
rect 50 108 60 109
<< ndcontact >>
rect 4 13 12 51
rect 30 12 38 50
rect 46 13 54 51
<< pdcontact >>
rect 4 149 12 187
rect 20 149 28 187
rect 36 116 44 184
rect 52 109 60 187
<< psubstratepcontact >>
rect -4 -4 4 4
rect 28 -4 36 4
<< nsubstratencontact >>
rect -4 196 4 204
rect 28 196 36 204
<< polysilicon >>
rect 14 188 18 192
rect 30 188 34 192
rect 46 188 50 192
rect 14 146 18 148
rect 10 142 18 146
rect 10 82 14 142
rect 12 74 14 82
rect 30 78 34 148
rect 10 60 14 74
rect 32 74 34 78
rect 10 56 18 60
rect 14 52 18 56
rect 24 52 28 70
rect 46 66 50 108
rect 48 62 50 66
rect 40 52 44 58
rect 14 8 18 12
rect 24 8 28 12
rect 40 8 44 12
<< polycontact >>
rect 4 74 12 82
rect 24 70 32 78
rect 40 58 48 66
<< metal1 >>
rect -4 204 68 206
rect 4 196 28 204
rect 36 196 68 204
rect -4 194 68 196
rect 4 187 12 194
rect 4 148 12 149
rect 20 187 28 188
rect 20 148 28 149
rect 22 106 28 148
rect 36 184 44 194
rect 36 112 44 116
rect 52 187 60 188
rect 52 108 60 109
rect 22 100 46 106
rect 20 86 28 94
rect 4 66 12 74
rect 22 78 28 86
rect 22 72 24 78
rect 40 66 46 100
rect 54 94 60 108
rect 52 86 60 94
rect 18 60 40 64
rect 6 58 40 60
rect 6 54 24 58
rect 6 52 12 54
rect 54 52 60 86
rect 4 51 12 52
rect 46 51 60 52
rect 4 12 12 13
rect 54 42 60 51
rect 46 12 54 13
rect 30 6 38 12
rect -4 4 68 6
rect 4 -4 28 4
rect 36 -4 68 4
rect -4 -6 68 -4
<< m1p >>
rect 20 86 28 94
rect 52 86 60 94
rect 4 66 12 74
<< labels >>
rlabel metal1 8 200 8 200 4 vdd
rlabel metal1 8 0 8 0 4 gnd
rlabel metal1 8 70 8 70 4 A
rlabel metal1 24 90 24 90 4 B
rlabel metal1 56 90 56 90 4 Y
<< end >>
