magic
tech scmos
magscale 1 2
timestamp 1600036665
<< checkpaint >>
rect -76 -66 428 270
<< nwell >>
rect -16 136 368 210
<< ntransistor >>
rect 16 12 20 52
rect 28 12 32 52
rect 48 12 52 52
rect 60 12 64 52
rect 94 12 98 32
rect 110 12 114 32
rect 126 12 130 32
rect 158 12 162 32
rect 174 12 178 32
rect 206 12 210 32
rect 222 12 226 32
rect 256 12 260 52
rect 268 12 272 52
rect 288 12 292 52
rect 300 12 304 52
rect 334 12 338 32
<< ptransistor >>
rect 14 148 18 188
rect 30 148 34 188
rect 46 148 50 188
rect 62 148 66 188
rect 94 168 98 188
rect 110 168 114 188
rect 126 148 130 188
rect 158 148 162 188
rect 174 148 178 188
rect 206 168 210 188
rect 222 168 226 188
rect 254 148 258 188
rect 270 148 274 188
rect 286 148 290 188
rect 302 148 306 188
rect 334 148 338 188
<< ndiffusion >>
rect 4 51 16 52
rect 12 13 16 51
rect 4 12 16 13
rect 20 12 28 52
rect 32 51 48 52
rect 32 13 36 51
rect 44 13 48 51
rect 32 12 48 13
rect 52 12 60 52
rect 64 51 76 52
rect 64 13 68 51
rect 244 51 256 52
rect 64 12 76 13
rect 84 31 94 32
rect 92 13 94 31
rect 84 12 94 13
rect 98 31 110 32
rect 98 13 100 31
rect 108 13 110 31
rect 98 12 110 13
rect 114 31 126 32
rect 114 13 116 31
rect 124 13 126 31
rect 114 12 126 13
rect 130 31 140 32
rect 130 13 132 31
rect 130 12 140 13
rect 148 31 158 32
rect 156 13 158 31
rect 148 12 158 13
rect 162 31 174 32
rect 162 13 164 31
rect 172 13 174 31
rect 162 12 174 13
rect 178 31 188 32
rect 178 13 180 31
rect 178 12 188 13
rect 196 31 206 32
rect 204 13 206 31
rect 196 12 206 13
rect 210 31 222 32
rect 210 13 212 31
rect 220 13 222 31
rect 210 12 222 13
rect 226 31 236 32
rect 226 13 228 31
rect 226 12 236 13
rect 252 13 256 51
rect 244 12 256 13
rect 260 12 268 52
rect 272 51 288 52
rect 272 13 276 51
rect 284 13 288 51
rect 272 12 288 13
rect 292 12 300 52
rect 304 51 316 52
rect 304 13 308 51
rect 304 12 316 13
rect 324 31 334 32
rect 332 13 334 31
rect 324 12 334 13
rect 338 31 348 32
rect 338 13 340 31
rect 338 12 348 13
<< pdiffusion >>
rect 4 187 14 188
rect 12 149 14 187
rect 4 148 14 149
rect 18 187 30 188
rect 18 149 20 187
rect 28 149 30 187
rect 18 148 30 149
rect 34 187 46 188
rect 34 149 36 187
rect 44 149 46 187
rect 34 148 46 149
rect 50 187 62 188
rect 50 149 52 187
rect 60 149 62 187
rect 50 148 62 149
rect 66 187 76 188
rect 66 149 68 187
rect 84 187 94 188
rect 92 169 94 187
rect 84 168 94 169
rect 98 187 110 188
rect 98 169 100 187
rect 108 169 110 187
rect 98 168 110 169
rect 114 187 126 188
rect 114 168 116 187
rect 66 148 76 149
rect 124 149 126 187
rect 116 148 126 149
rect 130 187 140 188
rect 130 149 132 187
rect 130 148 140 149
rect 148 187 158 188
rect 156 149 158 187
rect 148 148 158 149
rect 162 187 174 188
rect 162 149 164 187
rect 172 149 174 187
rect 162 148 174 149
rect 178 187 188 188
rect 178 149 180 187
rect 196 187 206 188
rect 204 169 206 187
rect 196 168 206 169
rect 210 187 222 188
rect 210 169 212 187
rect 220 169 222 187
rect 210 168 222 169
rect 226 187 236 188
rect 226 169 228 187
rect 226 168 236 169
rect 244 187 254 188
rect 178 148 188 149
rect 252 149 254 187
rect 244 148 254 149
rect 258 187 270 188
rect 258 149 260 187
rect 268 149 270 187
rect 258 148 270 149
rect 274 187 286 188
rect 274 149 276 187
rect 284 149 286 187
rect 274 148 286 149
rect 290 187 302 188
rect 290 149 292 187
rect 300 149 302 187
rect 290 148 302 149
rect 306 187 316 188
rect 306 149 308 187
rect 306 148 316 149
rect 324 187 334 188
rect 332 149 334 187
rect 324 148 334 149
rect 338 187 348 188
rect 338 149 340 187
rect 338 148 348 149
<< ndcontact >>
rect 4 13 12 51
rect 36 13 44 51
rect 68 13 76 51
rect 84 13 92 31
rect 100 13 108 31
rect 116 13 124 31
rect 132 13 140 31
rect 148 13 156 31
rect 164 13 172 31
rect 180 13 188 31
rect 196 13 204 31
rect 212 13 220 31
rect 228 13 236 31
rect 244 13 252 51
rect 276 13 284 51
rect 308 13 316 51
rect 324 13 332 31
rect 340 13 348 31
<< pdcontact >>
rect 4 149 12 187
rect 20 149 28 187
rect 36 149 44 187
rect 52 149 60 187
rect 68 149 76 187
rect 84 169 92 187
rect 100 169 108 187
rect 116 149 124 187
rect 132 149 140 187
rect 148 149 156 187
rect 164 149 172 187
rect 180 149 188 187
rect 196 169 204 187
rect 212 169 220 187
rect 228 169 236 187
rect 244 149 252 187
rect 260 149 268 187
rect 276 149 284 187
rect 292 149 300 187
rect 308 149 316 187
rect 324 149 332 187
rect 340 149 348 187
<< psubstratepcontact >>
rect -4 -4 4 4
rect 28 -4 36 4
rect 60 -4 68 4
rect 92 -4 100 4
rect 124 -4 132 4
rect 156 -4 164 4
rect 188 -4 196 4
rect 220 -4 228 4
rect 252 -4 260 4
rect 284 -4 292 4
<< nsubstratencontact >>
rect -4 196 4 204
rect 28 196 36 204
rect 60 196 68 204
rect 92 196 100 204
rect 124 196 132 204
rect 156 196 164 204
rect 188 196 196 204
rect 220 196 228 204
rect 252 196 260 204
rect 284 196 292 204
<< polysilicon >>
rect 14 188 18 192
rect 30 188 34 192
rect 46 188 50 192
rect 62 188 66 192
rect 94 188 98 192
rect 110 188 114 192
rect 126 188 130 192
rect 158 188 162 192
rect 174 188 178 192
rect 206 188 210 192
rect 222 188 226 192
rect 254 188 258 192
rect 270 188 274 192
rect 286 188 290 192
rect 302 188 306 192
rect 334 188 338 192
rect 14 146 18 148
rect 8 142 18 146
rect 8 96 12 142
rect 30 130 34 148
rect 28 122 34 130
rect 30 112 34 122
rect 46 128 50 148
rect 62 142 66 148
rect 94 146 98 168
rect 94 142 102 146
rect 62 138 70 142
rect 30 108 38 112
rect 8 88 18 96
rect 8 58 12 88
rect 34 66 38 108
rect 36 58 38 66
rect 46 58 50 120
rect 66 102 70 138
rect 62 98 70 102
rect 62 60 66 98
rect 98 84 102 142
rect 110 134 114 168
rect 206 166 210 168
rect 202 162 210 166
rect 126 146 130 148
rect 126 142 150 146
rect 110 126 130 134
rect 114 68 118 126
rect 146 118 150 142
rect 158 140 162 148
rect 174 146 178 148
rect 8 54 20 58
rect 16 52 20 54
rect 28 52 32 58
rect 46 54 52 58
rect 48 52 52 54
rect 60 56 66 60
rect 94 64 118 68
rect 126 114 150 118
rect 156 136 162 140
rect 168 142 178 146
rect 126 66 130 114
rect 156 84 160 136
rect 168 118 172 142
rect 202 134 206 162
rect 222 142 226 168
rect 188 126 206 134
rect 168 114 176 118
rect 60 52 64 56
rect 94 32 98 64
rect 126 58 132 66
rect 110 32 114 46
rect 126 32 130 58
rect 156 38 160 76
rect 172 54 176 114
rect 202 94 206 126
rect 200 90 206 94
rect 212 138 226 142
rect 192 62 194 70
rect 200 66 204 90
rect 212 82 220 138
rect 254 120 258 148
rect 270 146 274 148
rect 228 116 258 120
rect 266 142 274 146
rect 228 76 232 116
rect 266 108 270 142
rect 286 112 290 148
rect 258 104 270 108
rect 276 108 290 112
rect 302 108 306 148
rect 258 92 262 104
rect 252 84 262 92
rect 276 84 280 108
rect 228 72 240 76
rect 200 62 230 66
rect 190 54 194 62
rect 190 50 210 54
rect 156 34 162 38
rect 158 32 162 34
rect 174 32 178 46
rect 206 32 210 50
rect 226 38 230 62
rect 236 58 240 72
rect 258 68 262 84
rect 278 76 280 84
rect 276 68 280 76
rect 288 100 298 102
rect 288 98 306 100
rect 288 68 292 98
rect 334 84 338 148
rect 308 76 338 84
rect 258 64 270 68
rect 276 64 282 68
rect 288 64 304 68
rect 266 58 270 64
rect 278 58 282 64
rect 236 54 260 58
rect 266 54 272 58
rect 278 54 292 58
rect 256 52 260 54
rect 268 52 272 54
rect 288 52 292 54
rect 300 52 304 64
rect 222 34 230 38
rect 222 32 226 34
rect 334 32 338 76
rect 16 8 20 12
rect 28 8 32 12
rect 48 8 52 12
rect 60 8 64 12
rect 94 8 98 12
rect 110 8 114 12
rect 126 8 130 12
rect 158 8 162 12
rect 174 8 178 12
rect 206 8 210 12
rect 222 8 226 12
rect 256 8 260 12
rect 268 8 272 12
rect 288 8 292 12
rect 300 8 304 12
rect 334 8 338 12
<< polycontact >>
rect 20 122 28 130
rect 46 120 54 128
rect 18 88 26 96
rect 28 58 36 66
rect 70 102 78 110
rect 130 126 138 134
rect 98 76 106 84
rect 180 126 188 134
rect 156 76 164 84
rect 132 58 140 66
rect 110 46 118 54
rect 148 46 156 54
rect 184 62 192 70
rect 246 134 254 142
rect 212 74 220 82
rect 278 126 286 134
rect 244 84 252 92
rect 172 46 180 54
rect 210 46 218 54
rect 270 76 278 84
rect 298 100 306 108
rect 300 76 308 84
<< metal1 >>
rect -4 204 356 206
rect 4 196 28 204
rect 36 196 60 204
rect 68 196 92 204
rect 100 196 124 204
rect 132 196 156 204
rect 164 196 188 204
rect 196 196 220 204
rect 228 196 252 204
rect 260 196 284 204
rect 292 196 356 204
rect -4 194 356 196
rect 4 187 12 194
rect 20 187 28 188
rect 4 148 12 149
rect 18 149 20 154
rect 18 148 28 149
rect 36 187 44 194
rect 36 148 44 149
rect 52 187 60 188
rect 18 142 24 148
rect 52 142 60 149
rect 68 187 76 194
rect 84 187 92 188
rect 84 168 92 169
rect 100 187 108 188
rect 100 168 108 169
rect 116 187 124 188
rect 68 148 76 149
rect 116 148 124 149
rect 132 187 140 194
rect 132 148 140 149
rect 148 187 156 188
rect 148 148 156 149
rect 164 187 172 194
rect 164 148 172 149
rect 180 187 188 188
rect 196 187 204 188
rect 196 168 204 169
rect 212 187 220 188
rect 212 168 220 169
rect 228 187 236 188
rect 228 168 236 169
rect 244 187 252 194
rect 180 148 188 149
rect 244 148 252 149
rect 260 187 268 188
rect 4 136 24 142
rect 4 80 12 136
rect 30 134 72 142
rect 180 134 188 140
rect 220 134 246 142
rect 260 134 268 149
rect 276 187 284 194
rect 276 148 284 149
rect 292 187 300 188
rect 292 142 300 149
rect 308 187 316 194
rect 308 148 316 149
rect 324 187 332 188
rect 292 136 318 142
rect 30 130 36 134
rect 28 122 36 130
rect 66 128 124 134
rect 54 122 60 128
rect 54 116 100 122
rect 118 120 124 128
rect 138 126 148 134
rect 260 126 278 134
rect 118 114 196 120
rect 312 120 318 136
rect 236 114 318 120
rect 36 108 44 114
rect 36 102 70 108
rect 78 102 298 108
rect 312 96 318 114
rect 324 110 332 149
rect 340 187 348 194
rect 340 148 348 149
rect 324 102 334 110
rect 26 92 252 96
rect 26 90 244 92
rect 68 86 76 90
rect 312 90 320 96
rect 4 72 84 80
rect 106 76 118 84
rect 164 76 180 84
rect 4 51 12 72
rect 36 58 58 66
rect 50 52 58 58
rect 110 54 118 76
rect 132 66 140 74
rect 156 62 184 68
rect 212 54 220 74
rect 278 76 300 84
rect 270 64 278 76
rect 314 70 320 90
rect 4 12 12 13
rect 36 51 44 52
rect 50 51 76 52
rect 50 44 68 51
rect 36 6 44 13
rect 118 46 148 52
rect 164 46 172 54
rect 218 46 220 54
rect 260 58 278 64
rect 308 64 320 70
rect 260 52 268 58
rect 244 51 268 52
rect 68 12 76 13
rect 84 31 92 32
rect 84 12 92 13
rect 100 31 108 32
rect 100 12 108 13
rect 116 31 124 32
rect 116 12 124 13
rect 132 31 140 32
rect 132 6 140 13
rect 148 31 156 32
rect 148 12 156 13
rect 164 31 172 32
rect 164 6 172 13
rect 180 31 188 32
rect 180 12 188 13
rect 196 31 204 32
rect 196 12 204 13
rect 212 31 220 32
rect 212 12 220 13
rect 228 31 236 32
rect 228 12 236 13
rect 252 44 268 51
rect 276 51 284 52
rect 244 12 252 13
rect 276 6 284 13
rect 308 51 316 64
rect 326 58 334 102
rect 308 12 316 13
rect 324 50 334 58
rect 324 31 332 50
rect 324 12 332 13
rect 340 31 348 32
rect 340 6 348 13
rect -4 4 356 6
rect 4 -4 28 4
rect 36 -4 60 4
rect 68 -4 92 4
rect 100 -4 124 4
rect 132 -4 156 4
rect 164 -4 188 4
rect 196 -4 220 4
rect 228 -4 252 4
rect 260 -4 284 4
rect 292 -4 356 4
rect -4 -6 356 -4
<< m2contact >>
rect 84 160 92 168
rect 100 160 108 168
rect 196 160 204 168
rect 212 160 220 168
rect 228 160 236 168
rect 116 140 124 148
rect 148 140 156 148
rect 180 140 188 148
rect 212 134 220 142
rect 100 114 108 122
rect 148 126 156 134
rect 196 114 204 122
rect 228 114 236 122
rect 84 72 92 80
rect 180 76 188 84
rect 148 60 156 68
rect 84 32 92 40
rect 100 32 108 40
rect 116 32 124 40
rect 148 32 156 40
rect 180 32 188 40
rect 196 32 204 40
rect 212 32 220 40
rect 228 32 236 40
<< metal2 >>
rect 84 80 92 160
rect 84 40 92 72
rect 100 122 108 160
rect 100 40 108 114
rect 116 40 124 140
rect 148 134 156 140
rect 148 68 156 126
rect 148 40 156 60
rect 180 84 188 140
rect 180 40 188 76
rect 196 122 204 160
rect 196 40 204 114
rect 212 142 220 160
rect 212 40 220 134
rect 228 122 236 160
rect 228 40 236 114
<< m1p >>
rect 324 126 332 134
rect 36 106 44 114
rect 68 86 76 94
rect 132 66 140 74
rect 164 46 172 54
<< labels >>
rlabel metal1 8 0 8 0 4 gnd
rlabel metal1 8 200 8 200 4 vdd
rlabel metal1 136 70 136 70 4 D
rlabel metal1 40 110 40 110 4 S
rlabel metal1 72 90 72 90 4 R
rlabel metal1 328 130 328 130 4 Q
rlabel metal1 168 50 168 50 4 CLK
<< end >>
