magic
tech scmos
magscale 1 2
timestamp 1600036665
<< checkpaint >>
rect -76 -66 188 270
<< nwell >>
rect -16 96 128 210
<< ntransistor >>
rect 14 12 18 52
rect 32 12 36 52
rect 42 12 46 52
rect 66 12 70 52
rect 76 12 80 52
rect 94 12 98 52
<< ptransistor >>
rect 14 108 18 188
rect 32 108 36 188
rect 42 108 46 188
rect 66 108 70 188
rect 76 108 80 188
rect 94 108 98 188
<< ndiffusion >>
rect 4 51 14 52
rect 12 13 14 51
rect 4 12 14 13
rect 18 43 32 52
rect 18 15 21 43
rect 29 15 32 43
rect 18 12 32 15
rect 36 12 42 52
rect 46 44 66 52
rect 46 16 52 44
rect 60 16 66 44
rect 46 12 66 16
rect 70 12 76 52
rect 80 43 94 52
rect 80 15 83 43
rect 91 15 94 43
rect 80 12 94 15
rect 98 51 108 52
rect 98 13 100 51
rect 98 12 108 13
<< pdiffusion >>
rect 4 187 14 188
rect 12 109 14 187
rect 4 108 14 109
rect 18 184 32 188
rect 18 126 21 184
rect 29 126 32 184
rect 18 108 32 126
rect 36 108 42 188
rect 46 187 66 188
rect 46 109 52 187
rect 60 109 66 187
rect 46 108 66 109
rect 70 108 76 188
rect 80 184 94 188
rect 80 126 83 184
rect 91 126 94 184
rect 80 108 94 126
rect 98 187 108 188
rect 98 109 100 187
rect 98 108 108 109
<< ndcontact >>
rect 4 13 12 51
rect 21 15 29 43
rect 52 16 60 44
rect 83 15 91 43
rect 100 13 108 51
<< pdcontact >>
rect 4 109 12 187
rect 21 126 29 184
rect 52 109 60 187
rect 83 126 91 184
rect 100 109 108 187
<< psubstratepcontact >>
rect -4 -4 4 4
rect 28 -4 36 4
rect 60 -4 68 4
rect 92 -4 100 4
<< nsubstratencontact >>
rect -4 196 4 204
rect 28 196 36 204
rect 60 196 68 204
rect 92 196 100 204
<< polysilicon >>
rect 14 188 18 192
rect 32 188 36 192
rect 42 188 46 192
rect 66 188 70 192
rect 76 188 80 192
rect 94 188 98 192
rect 14 104 18 108
rect 32 106 36 108
rect 12 100 18 104
rect 28 102 36 106
rect 12 74 16 100
rect 28 90 32 102
rect 42 94 46 108
rect 14 52 18 66
rect 28 58 32 82
rect 50 74 54 94
rect 66 84 70 108
rect 76 106 80 108
rect 94 106 98 108
rect 76 102 98 106
rect 66 80 76 84
rect 72 74 76 80
rect 94 74 98 102
rect 50 70 64 74
rect 28 54 36 58
rect 32 52 36 54
rect 42 54 44 58
rect 60 58 64 70
rect 94 58 98 66
rect 60 54 70 58
rect 42 52 46 54
rect 66 52 70 54
rect 76 54 98 58
rect 76 52 80 54
rect 94 52 98 54
rect 14 8 18 12
rect 32 8 36 12
rect 42 8 46 12
rect 66 8 70 12
rect 76 8 80 12
rect 94 8 98 12
<< polycontact >>
rect 46 94 54 102
rect 24 82 32 90
rect 12 66 20 74
rect 44 54 52 62
rect 72 66 80 74
rect 92 66 100 74
<< metal1 >>
rect -4 204 116 206
rect 4 196 28 204
rect 36 196 60 204
rect 68 196 92 204
rect 100 196 116 204
rect -4 194 116 196
rect 22 188 30 194
rect 4 187 12 188
rect 20 184 30 188
rect 20 126 21 184
rect 29 126 30 184
rect 20 122 30 126
rect 48 187 64 188
rect 12 109 18 114
rect 4 108 18 109
rect 48 109 52 187
rect 60 114 64 187
rect 82 184 92 194
rect 82 126 83 184
rect 91 126 92 184
rect 82 122 92 126
rect 100 187 108 188
rect 60 109 68 114
rect 48 108 68 109
rect 92 109 100 114
rect 92 108 108 109
rect 20 102 26 108
rect 20 96 46 102
rect 62 94 68 108
rect 62 88 76 94
rect 32 82 50 88
rect 44 76 50 82
rect 58 86 76 88
rect 58 82 68 86
rect 4 66 12 74
rect 20 66 38 72
rect 32 62 38 66
rect 4 52 18 58
rect 32 56 36 62
rect 4 51 12 52
rect 58 48 64 82
rect 100 66 108 74
rect 72 62 78 66
rect 92 52 108 58
rect 4 12 12 13
rect 20 43 30 46
rect 20 15 21 43
rect 29 15 30 43
rect 20 12 30 15
rect 48 44 64 48
rect 100 51 108 52
rect 48 16 52 44
rect 60 16 64 44
rect 48 12 64 16
rect 82 43 92 46
rect 82 15 83 43
rect 91 15 92 43
rect 22 6 30 12
rect 82 6 92 15
rect 100 12 108 13
rect -4 4 116 6
rect 4 -4 28 4
rect 36 -4 60 4
rect 68 -4 92 4
rect 100 -4 116 4
rect -4 -6 116 -4
<< m2contact >>
rect 18 108 26 116
rect 84 108 92 116
rect 44 68 52 76
rect 18 52 26 60
rect 36 54 44 62
rect 70 54 78 62
rect 84 52 92 60
<< metal2 >>
rect 18 60 24 108
rect 86 74 92 108
rect 52 68 92 74
rect 44 54 70 60
rect 86 60 92 68
<< m1p >>
rect 68 86 76 94
rect 4 66 12 74
rect 100 66 108 74
<< labels >>
rlabel metal1 8 70 8 70 4 A
rlabel metal1 104 70 104 70 4 B
rlabel metal1 8 0 8 0 4 gnd
rlabel metal1 8 200 8 200 4 vdd
rlabel metal1 72 90 72 90 4 Y
<< end >>
